// TODO: implement this part

module ControlUnit (
  input [3:0] op_code,
  input [1:0] mode,
  input s_in,
  output s, b, exe_cmd, mem_w_en, mem_r_en, wb_en
  );

endmodule // ControlUnit
